LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY dataMem IS

	PORT(
		CLK : IN STD_LOGIC;
		MEMWR  : IN STD_LOGIC;
		RST : IN STD_LOGIC;
		-- 1kB
		ADDRESS : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		DATAIN  : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		M0 	: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		M1	: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		DATAOUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));

END ENTITY dataMem;


ARCHITECTURE dataMemArch OF dataMem IS
	
	TYPE RAM_TYPE IS ARRAY(0 TO 1023) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL DATAMEMORY : RAM_TYPE;
	SIGNAL M0ADD : std_logic_vector(9 downto 0);
	SIGNAL M1ADD : std_logic_vector(9 downto 0);
	BEGIN
		M0ADD <= "0000000000";
		M1ADD <= "0000000001";

		PROCESS(CLK, RST) IS -- WRITE ON RISING EDGE (Sync.)
			BEGIN
				IF RST = '1' THEN
					DATAMEMORY <= (others => (others => '0'));
				ELSIF RISING_EDGE(CLK) THEN
					IF MEMWR = '1' THEN
						DATAMEMORY (TO_INTEGER(UNSIGNED(ADDRESS))) <= DATAIN;
					END IF;
				END IF;
		END PROCESS;
		
		DATAOUT <= DATAMEMORY (TO_INTEGER(UNSIGNED(ADDRESS))); -- Async.
		M0 <= DATAMEMORY (TO_INTEGER(UNSIGNED(M0ADD)));
		M1 <= DATAMEMORY (TO_INTEGER(UNSIGNED(M1ADD)));
END dataMemArch;