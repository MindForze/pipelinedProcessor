LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY instMem IS
	PORT(
		--1KB ADD.SPACE BUT PC IS 16 BITS
		ADDRESS : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		INSTOUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END ENTITY instMem;

ARCHITECTURE instMemArch OF instMem IS
	
	TYPE RAM_TYPE IS ARRAY(0 TO 1023) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL MEMORY : RAM_TYPE;

	BEGIN
	INSTOUT <= MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)));


END instMemArch;
